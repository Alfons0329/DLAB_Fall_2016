`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:13:08 12/31/2016 
// Design Name: 
// Module Name:    state 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module state(
    output reg stateleft,
    output reg statedown,
    output reg stateup,
	output reg statew,
	output reg states,
	output reg stated,
    input clk,
    input rst,
    input [9:0] Data
    );
    
always@(posedge clk, posedge rst) begin
    if(rst) stateleft <= 0;
    else begin
        case(Data)
        {2'b01,8'h6B}: stateleft <= 1;
        {2'b11,8'h6B}: stateleft <= 0;
        default: stateleft <= stateleft;
        endcase
    end
end

always@(posedge clk, posedge rst) begin
    if(rst) stateup <= 0;
    else begin
        case(Data)
        {2'b01,8'h75}: stateup <= 1;
        {2'b11,8'h75}: stateup <= 0;
        default: stateup <= stateup;
        endcase
    end
end

always@(posedge clk, posedge rst) begin
    if(rst) statedown <= 0;
    else begin
        case(Data)
        {2'b01,8'h72}: statedown <= 1;
        {2'b11,8'h72}: statedown <= 0;
        default: statedown <= statedown;
        endcase
    end
end

///////WSD

//W
always@(posedge clk, posedge rst) begin
    if(rst) statew <= 0;
    else begin
        case(Data)
        {2'b00,8'h1D}: statew <= 1;
        {2'b10,8'h1D}: statew <= 0;
        default: statew <= statew;
        endcase
    end
end
//S
always@(posedge clk, posedge rst) begin
    if(rst) states <= 0;
    else begin
        case(Data)
        {2'b00,8'h1B}: states <= 1;
        {2'b10,8'h1B}: states <= 0;
        default: states <= states;
        endcase
    end
end
//D
always@(posedge clk, posedge rst) begin
    if(rst) stated <= 0;
    else begin
        case(Data)
        {2'b00,8'h23}: stated <= 1;
        {2'b10,8'h23}: stated <= 0;
        default: stated <= stated;
        endcase
    end
end


endmodule
